// niosmp.v

// Generated using ACDS version 14.0 200 at 2015.12.06.20:50:11

`timescale 1 ps / 1 ps
module niosmp (
		input  wire       clk_clk,          //       clk.clk
		input  wire       reset_reset_n,    //     reset.reset_n
		output wire [7:0] leds_export,      //      leds.export
		inout  wire [7:0] data_export,      //      data.export
		output wire [7:0] address_export,   //   address.export
		output wire       rnw_export,       //       rnw.export
		output wire       noe_export,       //       noe.export
		input  wire [7:0] mpdatain_export,  //  mpdatain.export
		input  wire       chrec_export,     //     chrec.export
		output wire [7:0] mpdataout_export, // mpdataout.export
		output wire       asoe_export,      //      asoe.export
		input  wire       sent_export,      //      sent.export
		output wire       load_export,      //      load.export
		input  wire       testin_export     //    testin.export
	);

	wire         nios2_processor_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [19:0] nios2_processor_instruction_master_address;                      // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                         // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire  [31:0] nios2_processor_instruction_master_readdata;                     // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_processor_instruction_master_readdatavalid -> nios2_processor:i_readdatavalid
	wire         nios2_processor_data_master_waitrequest;                         // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire  [31:0] nios2_processor_data_master_writedata;                           // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [19:0] nios2_processor_data_master_address;                             // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire         nios2_processor_data_master_write;                               // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire         nios2_processor_data_master_read;                                // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire  [31:0] nios2_processor_data_master_readdata;                            // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_debugaccess;                         // nios2_processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire         nios2_processor_data_master_readdatavalid;                       // mm_interconnect_0:nios2_processor_data_master_readdatavalid -> nios2_processor:d_readdatavalid
	wire   [3:0] nios2_processor_data_master_byteenable;                          // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest; // nios2_processor:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_processor_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_processor_jtag_debug_module_writedata -> nios2_processor:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_processor_jtag_debug_module_address;     // mm_interconnect_0:nios2_processor_jtag_debug_module_address -> nios2_processor:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_write;       // mm_interconnect_0:nios2_processor_jtag_debug_module_write -> nios2_processor:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_read;        // mm_interconnect_0:nios2_processor_jtag_debug_module_read -> nios2_processor:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_readdata;    // nios2_processor:jtag_debug_module_readdata -> mm_interconnect_0:nios2_processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_processor_jtag_debug_module_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_processor_jtag_debug_module_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                    // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                      // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                   // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;                        // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;                        // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                     // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                   // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                             // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                               // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_chipselect;                            // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire         mm_interconnect_0_leds_s1_write;                                 // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                              // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_data_s1_writedata;                             // mm_interconnect_0:data_s1_writedata -> data:writedata
	wire   [1:0] mm_interconnect_0_data_s1_address;                               // mm_interconnect_0:data_s1_address -> data:address
	wire         mm_interconnect_0_data_s1_chipselect;                            // mm_interconnect_0:data_s1_chipselect -> data:chipselect
	wire         mm_interconnect_0_data_s1_write;                                 // mm_interconnect_0:data_s1_write -> data:write_n
	wire  [31:0] mm_interconnect_0_data_s1_readdata;                              // data:readdata -> mm_interconnect_0:data_s1_readdata
	wire  [31:0] mm_interconnect_0_address_s1_writedata;                          // mm_interconnect_0:address_s1_writedata -> address:writedata
	wire   [1:0] mm_interconnect_0_address_s1_address;                            // mm_interconnect_0:address_s1_address -> address:address
	wire         mm_interconnect_0_address_s1_chipselect;                         // mm_interconnect_0:address_s1_chipselect -> address:chipselect
	wire         mm_interconnect_0_address_s1_write;                              // mm_interconnect_0:address_s1_write -> address:write_n
	wire  [31:0] mm_interconnect_0_address_s1_readdata;                           // address:readdata -> mm_interconnect_0:address_s1_readdata
	wire  [31:0] mm_interconnect_0_rnw_s1_writedata;                              // mm_interconnect_0:rnw_s1_writedata -> rnw:writedata
	wire   [1:0] mm_interconnect_0_rnw_s1_address;                                // mm_interconnect_0:rnw_s1_address -> rnw:address
	wire         mm_interconnect_0_rnw_s1_chipselect;                             // mm_interconnect_0:rnw_s1_chipselect -> rnw:chipselect
	wire         mm_interconnect_0_rnw_s1_write;                                  // mm_interconnect_0:rnw_s1_write -> rnw:write_n
	wire  [31:0] mm_interconnect_0_rnw_s1_readdata;                               // rnw:readdata -> mm_interconnect_0:rnw_s1_readdata
	wire  [31:0] mm_interconnect_0_noe_s1_writedata;                              // mm_interconnect_0:noe_s1_writedata -> noe:writedata
	wire   [1:0] mm_interconnect_0_noe_s1_address;                                // mm_interconnect_0:noe_s1_address -> noe:address
	wire         mm_interconnect_0_noe_s1_chipselect;                             // mm_interconnect_0:noe_s1_chipselect -> noe:chipselect
	wire         mm_interconnect_0_noe_s1_write;                                  // mm_interconnect_0:noe_s1_write -> noe:write_n
	wire  [31:0] mm_interconnect_0_noe_s1_readdata;                               // noe:readdata -> mm_interconnect_0:noe_s1_readdata
	wire   [1:0] mm_interconnect_0_mpdatain_s1_address;                           // mm_interconnect_0:mpdatain_s1_address -> mpdatain:address
	wire  [31:0] mm_interconnect_0_mpdatain_s1_readdata;                          // mpdatain:readdata -> mm_interconnect_0:mpdatain_s1_readdata
	wire   [1:0] mm_interconnect_0_chrec_s1_address;                              // mm_interconnect_0:chrec_s1_address -> chrec:address
	wire  [31:0] mm_interconnect_0_chrec_s1_readdata;                             // chrec:readdata -> mm_interconnect_0:chrec_s1_readdata
	wire  [31:0] mm_interconnect_0_mpdataout_s1_writedata;                        // mm_interconnect_0:mpdataout_s1_writedata -> mpdataout:writedata
	wire   [1:0] mm_interconnect_0_mpdataout_s1_address;                          // mm_interconnect_0:mpdataout_s1_address -> mpdataout:address
	wire         mm_interconnect_0_mpdataout_s1_chipselect;                       // mm_interconnect_0:mpdataout_s1_chipselect -> mpdataout:chipselect
	wire         mm_interconnect_0_mpdataout_s1_write;                            // mm_interconnect_0:mpdataout_s1_write -> mpdataout:write_n
	wire  [31:0] mm_interconnect_0_mpdataout_s1_readdata;                         // mpdataout:readdata -> mm_interconnect_0:mpdataout_s1_readdata
	wire  [31:0] mm_interconnect_0_asoe_s1_writedata;                             // mm_interconnect_0:asoe_s1_writedata -> asoe:writedata
	wire   [1:0] mm_interconnect_0_asoe_s1_address;                               // mm_interconnect_0:asoe_s1_address -> asoe:address
	wire         mm_interconnect_0_asoe_s1_chipselect;                            // mm_interconnect_0:asoe_s1_chipselect -> asoe:chipselect
	wire         mm_interconnect_0_asoe_s1_write;                                 // mm_interconnect_0:asoe_s1_write -> asoe:write_n
	wire  [31:0] mm_interconnect_0_asoe_s1_readdata;                              // asoe:readdata -> mm_interconnect_0:asoe_s1_readdata
	wire   [1:0] mm_interconnect_0_sent_s1_address;                               // mm_interconnect_0:sent_s1_address -> sent:address
	wire  [31:0] mm_interconnect_0_sent_s1_readdata;                              // sent:readdata -> mm_interconnect_0:sent_s1_readdata
	wire  [31:0] mm_interconnect_0_load_s1_writedata;                             // mm_interconnect_0:load_s1_writedata -> load:writedata
	wire   [1:0] mm_interconnect_0_load_s1_address;                               // mm_interconnect_0:load_s1_address -> load:address
	wire         mm_interconnect_0_load_s1_chipselect;                            // mm_interconnect_0:load_s1_chipselect -> load:chipselect
	wire         mm_interconnect_0_load_s1_write;                                 // mm_interconnect_0:load_s1_write -> load:write_n
	wire  [31:0] mm_interconnect_0_load_s1_readdata;                              // load:readdata -> mm_interconnect_0:load_s1_readdata
	wire   [1:0] mm_interconnect_0_testin_s1_address;                             // mm_interconnect_0:testin_s1_address -> testin:address
	wire  [31:0] mm_interconnect_0_testin_s1_readdata;                            // testin:readdata -> mm_interconnect_0:testin_s1_readdata
	wire         irq_mapper_receiver0_irq;                                        // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_processor_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:d_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [LEDs:reset_n, address:reset_n, asoe:reset_n, chrec:reset_n, data:reset_n, irq_mapper:reset, load:reset_n, mm_interconnect_0:nios2_processor_reset_n_reset_bridge_in_reset_reset, mpdatain:reset_n, mpdataout:reset_n, nios2_processor:reset_n, noe:reset_n, onchip_memory:reset, rnw:reset_n, rst_translator:in_reset, sent:reset_n, testin:reset_n]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_processor_jtag_debug_module_reset_reset;                   // nios2_processor:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset]

	niosmp_nios2_processor nios2_processor (
		.clk                                   (clk_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                              //                          .reset_req
		.d_address                             (nios2_processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                               //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_processor_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_processor_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                 // custom_instruction_master.readra
	);

	niosmp_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	niosmp_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	niosmp_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	niosmp_data data (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_s1_readdata),   //                    .readdata
		.bidir_port (data_export)                           // external_connection.export
	);

	niosmp_LEDs address (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_address_s1_readdata),   //                    .readdata
		.out_port   (address_export)                           // external_connection.export
	);

	niosmp_rnw rnw (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_rnw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rnw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rnw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rnw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rnw_s1_readdata),   //                    .readdata
		.out_port   (rnw_export)                           // external_connection.export
	);

	niosmp_rnw noe (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_noe_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_noe_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_noe_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_noe_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_noe_s1_readdata),   //                    .readdata
		.out_port   (noe_export)                           // external_connection.export
	);

	niosmp_mpdatain mpdatain (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_mpdatain_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_mpdatain_s1_readdata), //                    .readdata
		.in_port  (mpdatain_export)                         // external_connection.export
	);

	niosmp_chrec chrec (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_chrec_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_chrec_s1_readdata), //                    .readdata
		.in_port  (chrec_export)                         // external_connection.export
	);

	niosmp_LEDs mpdataout (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_mpdataout_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mpdataout_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mpdataout_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mpdataout_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mpdataout_s1_readdata),   //                    .readdata
		.out_port   (mpdataout_export)                           // external_connection.export
	);

	niosmp_rnw asoe (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_asoe_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_asoe_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_asoe_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_asoe_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_asoe_s1_readdata),   //                    .readdata
		.out_port   (asoe_export)                           // external_connection.export
	);

	niosmp_chrec sent (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_sent_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sent_s1_readdata), //                    .readdata
		.in_port  (sent_export)                         // external_connection.export
	);

	niosmp_rnw load (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_load_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_load_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_load_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_load_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_load_s1_readdata),   //                    .readdata
		.out_port   (load_export)                           // external_connection.export
	);

	niosmp_chrec testin (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_testin_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_testin_s1_readdata), //                    .readdata
		.in_port  (testin_export)                         // external_connection.export
	);

	niosmp_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                         //                                     clk_0_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                              //         jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // nios2_processor_reset_n_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address                 (nios2_processor_data_master_address),                             //                   nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest             (nios2_processor_data_master_waitrequest),                         //                                              .waitrequest
		.nios2_processor_data_master_byteenable              (nios2_processor_data_master_byteenable),                          //                                              .byteenable
		.nios2_processor_data_master_read                    (nios2_processor_data_master_read),                                //                                              .read
		.nios2_processor_data_master_readdata                (nios2_processor_data_master_readdata),                            //                                              .readdata
		.nios2_processor_data_master_readdatavalid           (nios2_processor_data_master_readdatavalid),                       //                                              .readdatavalid
		.nios2_processor_data_master_write                   (nios2_processor_data_master_write),                               //                                              .write
		.nios2_processor_data_master_writedata               (nios2_processor_data_master_writedata),                           //                                              .writedata
		.nios2_processor_data_master_debugaccess             (nios2_processor_data_master_debugaccess),                         //                                              .debugaccess
		.nios2_processor_instruction_master_address          (nios2_processor_instruction_master_address),                      //            nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest      (nios2_processor_instruction_master_waitrequest),                  //                                              .waitrequest
		.nios2_processor_instruction_master_read             (nios2_processor_instruction_master_read),                         //                                              .read
		.nios2_processor_instruction_master_readdata         (nios2_processor_instruction_master_readdata),                     //                                              .readdata
		.nios2_processor_instruction_master_readdatavalid    (nios2_processor_instruction_master_readdatavalid),                //                                              .readdatavalid
		.address_s1_address                                  (mm_interconnect_0_address_s1_address),                            //                                    address_s1.address
		.address_s1_write                                    (mm_interconnect_0_address_s1_write),                              //                                              .write
		.address_s1_readdata                                 (mm_interconnect_0_address_s1_readdata),                           //                                              .readdata
		.address_s1_writedata                                (mm_interconnect_0_address_s1_writedata),                          //                                              .writedata
		.address_s1_chipselect                               (mm_interconnect_0_address_s1_chipselect),                         //                                              .chipselect
		.asoe_s1_address                                     (mm_interconnect_0_asoe_s1_address),                               //                                       asoe_s1.address
		.asoe_s1_write                                       (mm_interconnect_0_asoe_s1_write),                                 //                                              .write
		.asoe_s1_readdata                                    (mm_interconnect_0_asoe_s1_readdata),                              //                                              .readdata
		.asoe_s1_writedata                                   (mm_interconnect_0_asoe_s1_writedata),                             //                                              .writedata
		.asoe_s1_chipselect                                  (mm_interconnect_0_asoe_s1_chipselect),                            //                                              .chipselect
		.chrec_s1_address                                    (mm_interconnect_0_chrec_s1_address),                              //                                      chrec_s1.address
		.chrec_s1_readdata                                   (mm_interconnect_0_chrec_s1_readdata),                             //                                              .readdata
		.data_s1_address                                     (mm_interconnect_0_data_s1_address),                               //                                       data_s1.address
		.data_s1_write                                       (mm_interconnect_0_data_s1_write),                                 //                                              .write
		.data_s1_readdata                                    (mm_interconnect_0_data_s1_readdata),                              //                                              .readdata
		.data_s1_writedata                                   (mm_interconnect_0_data_s1_writedata),                             //                                              .writedata
		.data_s1_chipselect                                  (mm_interconnect_0_data_s1_chipselect),                            //                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                              .chipselect
		.LEDs_s1_address                                     (mm_interconnect_0_leds_s1_address),                               //                                       LEDs_s1.address
		.LEDs_s1_write                                       (mm_interconnect_0_leds_s1_write),                                 //                                              .write
		.LEDs_s1_readdata                                    (mm_interconnect_0_leds_s1_readdata),                              //                                              .readdata
		.LEDs_s1_writedata                                   (mm_interconnect_0_leds_s1_writedata),                             //                                              .writedata
		.LEDs_s1_chipselect                                  (mm_interconnect_0_leds_s1_chipselect),                            //                                              .chipselect
		.load_s1_address                                     (mm_interconnect_0_load_s1_address),                               //                                       load_s1.address
		.load_s1_write                                       (mm_interconnect_0_load_s1_write),                                 //                                              .write
		.load_s1_readdata                                    (mm_interconnect_0_load_s1_readdata),                              //                                              .readdata
		.load_s1_writedata                                   (mm_interconnect_0_load_s1_writedata),                             //                                              .writedata
		.load_s1_chipselect                                  (mm_interconnect_0_load_s1_chipselect),                            //                                              .chipselect
		.mpdatain_s1_address                                 (mm_interconnect_0_mpdatain_s1_address),                           //                                   mpdatain_s1.address
		.mpdatain_s1_readdata                                (mm_interconnect_0_mpdatain_s1_readdata),                          //                                              .readdata
		.mpdataout_s1_address                                (mm_interconnect_0_mpdataout_s1_address),                          //                                  mpdataout_s1.address
		.mpdataout_s1_write                                  (mm_interconnect_0_mpdataout_s1_write),                            //                                              .write
		.mpdataout_s1_readdata                               (mm_interconnect_0_mpdataout_s1_readdata),                         //                                              .readdata
		.mpdataout_s1_writedata                              (mm_interconnect_0_mpdataout_s1_writedata),                        //                                              .writedata
		.mpdataout_s1_chipselect                             (mm_interconnect_0_mpdataout_s1_chipselect),                       //                                              .chipselect
		.nios2_processor_jtag_debug_module_address           (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //             nios2_processor_jtag_debug_module.address
		.nios2_processor_jtag_debug_module_write             (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                                              .write
		.nios2_processor_jtag_debug_module_read              (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                                              .read
		.nios2_processor_jtag_debug_module_readdata          (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                                              .readdata
		.nios2_processor_jtag_debug_module_writedata         (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                                              .writedata
		.nios2_processor_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                                              .byteenable
		.nios2_processor_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                                              .waitrequest
		.nios2_processor_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                                              .debugaccess
		.noe_s1_address                                      (mm_interconnect_0_noe_s1_address),                                //                                        noe_s1.address
		.noe_s1_write                                        (mm_interconnect_0_noe_s1_write),                                  //                                              .write
		.noe_s1_readdata                                     (mm_interconnect_0_noe_s1_readdata),                               //                                              .readdata
		.noe_s1_writedata                                    (mm_interconnect_0_noe_s1_writedata),                              //                                              .writedata
		.noe_s1_chipselect                                   (mm_interconnect_0_noe_s1_chipselect),                             //                                              .chipselect
		.onchip_memory_s1_address                            (mm_interconnect_0_onchip_memory_s1_address),                      //                              onchip_memory_s1.address
		.onchip_memory_s1_write                              (mm_interconnect_0_onchip_memory_s1_write),                        //                                              .write
		.onchip_memory_s1_readdata                           (mm_interconnect_0_onchip_memory_s1_readdata),                     //                                              .readdata
		.onchip_memory_s1_writedata                          (mm_interconnect_0_onchip_memory_s1_writedata),                    //                                              .writedata
		.onchip_memory_s1_byteenable                         (mm_interconnect_0_onchip_memory_s1_byteenable),                   //                                              .byteenable
		.onchip_memory_s1_chipselect                         (mm_interconnect_0_onchip_memory_s1_chipselect),                   //                                              .chipselect
		.onchip_memory_s1_clken                              (mm_interconnect_0_onchip_memory_s1_clken),                        //                                              .clken
		.rnw_s1_address                                      (mm_interconnect_0_rnw_s1_address),                                //                                        rnw_s1.address
		.rnw_s1_write                                        (mm_interconnect_0_rnw_s1_write),                                  //                                              .write
		.rnw_s1_readdata                                     (mm_interconnect_0_rnw_s1_readdata),                               //                                              .readdata
		.rnw_s1_writedata                                    (mm_interconnect_0_rnw_s1_writedata),                              //                                              .writedata
		.rnw_s1_chipselect                                   (mm_interconnect_0_rnw_s1_chipselect),                             //                                              .chipselect
		.sent_s1_address                                     (mm_interconnect_0_sent_s1_address),                               //                                       sent_s1.address
		.sent_s1_readdata                                    (mm_interconnect_0_sent_s1_readdata),                              //                                              .readdata
		.testin_s1_address                                   (mm_interconnect_0_testin_s1_address),                             //                                     testin_s1.address
		.testin_s1_readdata                                  (mm_interconnect_0_testin_s1_readdata)                             //                                              .readdata
	);

	niosmp_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                                // reset_in0.reset
		.reset_in1      (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),            //          .reset_req
		.reset_req_in0  (1'b0),                                          // (terminated)
		.reset_req_in1  (1'b0),                                          // (terminated)
		.reset_in2      (1'b0),                                          // (terminated)
		.reset_req_in2  (1'b0),                                          // (terminated)
		.reset_in3      (1'b0),                                          // (terminated)
		.reset_req_in3  (1'b0),                                          // (terminated)
		.reset_in4      (1'b0),                                          // (terminated)
		.reset_req_in4  (1'b0),                                          // (terminated)
		.reset_in5      (1'b0),                                          // (terminated)
		.reset_req_in5  (1'b0),                                          // (terminated)
		.reset_in6      (1'b0),                                          // (terminated)
		.reset_req_in6  (1'b0),                                          // (terminated)
		.reset_in7      (1'b0),                                          // (terminated)
		.reset_req_in7  (1'b0),                                          // (terminated)
		.reset_in8      (1'b0),                                          // (terminated)
		.reset_req_in8  (1'b0),                                          // (terminated)
		.reset_in9      (1'b0),                                          // (terminated)
		.reset_req_in9  (1'b0),                                          // (terminated)
		.reset_in10     (1'b0),                                          // (terminated)
		.reset_req_in10 (1'b0),                                          // (terminated)
		.reset_in11     (1'b0),                                          // (terminated)
		.reset_req_in11 (1'b0),                                          // (terminated)
		.reset_in12     (1'b0),                                          // (terminated)
		.reset_req_in12 (1'b0),                                          // (terminated)
		.reset_in13     (1'b0),                                          // (terminated)
		.reset_req_in13 (1'b0),                                          // (terminated)
		.reset_in14     (1'b0),                                          // (terminated)
		.reset_req_in14 (1'b0),                                          // (terminated)
		.reset_in15     (1'b0),                                          // (terminated)
		.reset_req_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
